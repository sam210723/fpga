module spdif (
  input CLK     // S/PDIF Clock
);

endmodule
