/*
 *  nco.v
 *  http://github.com/sam210723/fpga
 *
 *  Numerically Controlled Ocillator for a logic Phase-locked Loop.
 *
 */

module nco(
    input clk
);

    

endmodule
