module i2c_peripheral (
    inout           SDA,
    input           SCL,
    
    output  [7:0]   LED,
    output          OK
);

endmodule
