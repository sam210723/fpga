module i2c_controller (
    inout       SDA,
    output      SCL
);

    assign SDA = 0;
    assign SCL = 0;

endmodule
