module pma (
    input  clk,     // 250 MHz Ethernet Clock

);

    );

endmodule

