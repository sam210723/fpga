module spdif (
  input  clock    // S/PDIF Clock
);

endmodule
