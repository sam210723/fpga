module top(
    input       CLK_100MHz
);

endmodule
