/*
 *  nco.v
 *  http://github.com/sam210723/fpga
 *
 *  Numerically Controlled Oscillator for a logic Phase-locked Loop.
 *
 */

module nco(
    input clk
);

    

endmodule
